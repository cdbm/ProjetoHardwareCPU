module J5B( input wire [15:0] J20F, output wire [5:0] JFio);

assign JFio = J20F[5:0];

endmodule 